module simple_circuit(A2,B2,C2,Y);

output Y;

input A2,B2,C2;

wire w1,w2,w3;

assign w1= --------------------;
assign w2= --------------------;
assign w3= ------------------; 
assign Y=   -----------------;
 
endmodule
