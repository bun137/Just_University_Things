module not1( a,c );
--------------
-------------
-------------;
endmodule
