module xnor2( a,b,c);
input a,b;
output c;
assign c= ------------- ;
endmodule