module dfrl_16 (input wire  clk, reset, load, input wire [0:15] in, output wire [0:15] out);
  dfrl dfrl_0(clk, reset, load, in[0], out[0]);
  dfrl dfrl_1(--------------------------------);
  dfrl dfrl_2(--------------------------------);
  dfrl dfrl_3(--------------------------------);
  dfrl dfrl_4(--------------------------------);
  dfrl dfrl_5(--------------------------------);
  dfrl dfrl_6(--------------------------------);
  dfrl dfrl_7(--------------------------------);
  dfrl dfrl_8(-------------------------------);
  dfrl dfrl_9(----------------------);
  dfrl dfrl_10(----------------------);
  dfrl dfrl_11(----------------------);
  dfrl dfrl_12(----------------------);
  dfrl dfrl_13(----------------------);
  dfrl dfrl_14(----------------------);
  dfrl dfrl_15(----------------------);
endmodule

module mux2_16 (input wire [15:0] i0, i1, input wire j, output wire [15:0] o);
  mux2 mux2_0 (----------------------);
  mux2 mux2_1 (----------------------);
  mux2 mux2_2 (----------------------);
  mux2 mux2_3 (----------------------);
  mux2 mux2_4 (----------------------);
  mux2 mux2_5 (----------------------);
  mux2 mux2_6 (----------------------);
  mux2 mux2_7 (----------------------);
  mux2 mux2_8 (----------------------);
  mux2 mux2_9 (----------------------);
  mux2 mux2_10 (----------------------);
  mux2 mux2_11 (----------------------);
  mux2 mux2_12 (----------------------);
  mux2 mux2_13 (----------------------);
  mux2 mux2_14 (----------------------);
  mux2 mux2_15 (----------------------);
endmodule

module mux8_16 (input wire [0:15] i0, i1, i2, i3, i4, i5, i6, i7, input wire [0:2] j, output wire [0:15] o);
  mux8 mux8_0({i0[0], i1[0], i2[0], i3[0], i4[0], i5[0], i6[0], i7[0]}, j[0], j[1], j[2], o[0]);
  mux8 mux8_1(--------------------------------);
  mux8 mux8_2(--------------------------------);
  mux8 mux8_3(--------------------------------);
  mux8 mux8_4(--------------------------------);
  mux8 mux8_5(--------------------------------);
  mux8 mux8_6(--------------------------------);
  mux8 mux8_7(--------------------------------);
  mux8 mux8_8(--------------------------------);
  mux8 mux8_9(--------------------------------);
  mux8 mux8_10(-------------------------------);
  mux8 mux8_11(-------------------------------);
  mux8 mux8_12(-------------------------------);
  mux8 mux8_13(-------------------------------);
  mux8 mux8_14(-------------------------------);
  mux8 mux8_15(-------------------------------);
endmodule

module reg_file (input wire  clk, reset, wr, input wire [0:2] rd_addr_a, rd_addr_b, wr_addr, input wire [0:15] d_in, output wire [0:15] d_out_a, d_out_b);
  wire [0:7] load;  wire [0:15] dout_0, dout_1, dout_2, dout_3, dout_4, dout_5, dout_6, dout_7;

  dfrl_16 dfrl_16_0(clk, reset, load[0], d_in, dout_0);
  dfrl_16 dfrl_16_1(--------------------------------);
  dfrl_16 dfrl_16_2(--------------------------------);
  dfrl_16 dfrl_16_3(--------------------------------);
  dfrl_16 dfrl_16_4(--------------------------------);
  dfrl_16 dfrl_16_5(--------------------------------);
  dfrl_16 dfrl_16_6(------------------------------);
  dfrl_16 dfrl_16_7(--------------------------------);
  demux8 demux8_0(--------------------------------);
  mux8_16 mux8_16_9(----------------------);
  mux8_16 mux8_16_10(--------------------------------);
endmodule

module reg_alu (input wire clk, reset, sel, wr, input wire [1:0] op, input wire [2:0] rd_addr_a,
  rd_addr_b, wr_addr, input wire [15:0] d_in, output wire [15:0] d_out_a, d_out_b, output wire cout);
  wire [15:0] d_in_alu, d_in_reg; wire cout_0;
  alu alu_0 (--------------------------------);
  reg_file reg_file_0 (--------------------------------);
  mux2_16 mux2_16_0 (--------------------------------);
  dfr dfr_0 (--------------------------------);
endmodule
