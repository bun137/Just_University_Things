module simple_circuit(A,B,C,D,E);

output D,E;

input A,B,C;

wire w1;

and G1(------------);

not G2(------------);

or G3(------------);

endmodule
