module nor2( a,b,c);
-----------------
-----------------
----------------- ;
endmodule
